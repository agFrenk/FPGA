library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity encoder_rle_reset_tb is
end encoder_rle_reset_tb;

architecture testbench_architecture of encoder_rle_reset_tb is
    -- Constants
    constant WIDTH : natural := 64;
    
    -- Signals
    signal input_sig                : std_logic_vector(WIDTH-1 downto 0);
    signal clk_sig                  : std_logic := '0';
    signal reset_sig                : std_logic := '0';
    signal output_sig               : std_logic_vector((WIDTH*2)-1 downto 0);
    signal ready_sig                : std_logic;
    signal size_sig                 : integer;
    signal input_signal_ready_sig   : std_logic;



    -- Component declaration
    component encoder_rle
        generic (WIDTH : natural := 64);
        port (
            input_i                 : in std_logic_vector(WIDTH-1 downto 0);
            clk_i                   : in std_logic;
            reset_i                 : in std_logic;
            output_o                : out std_logic_vector((WIDTH*2)-1 downto 0);
            ready_o                 : out std_logic;
            input_signal_ready_i    : in std_logic;
            size_o                  : out integer
        );
    end component;

begin
    -- DUT instantiation
    uut: encoder_rle
    generic map (
        WIDTH => WIDTH
    )
    port map (
        input_i                 => input_sig,
        clk_i                   => clk_sig,
        reset_i                 => reset_sig,
        output_o                => output_sig,
        ready_o                 => ready_sig,
        input_signal_ready_i    => input_signal_ready_sig,
        size_o                  => size_sig
    );

    -- Clock generation process
    process
    begin
        while now < 1000 ns loop
            clk_sig <= '0';
            wait for 5 ns;
            clk_sig <= '1';
            wait for 5 ns;
        end loop;
        wait;
    end process;

    -- Stimulus process
    process
    begin
        -- Provide test vector
        input_signal_ready_sig <= '1';
        input_sig <= "1111111110101010101010101111000011000000101110101111010111110101";
        wait for 10 ns;
        input_signal_ready_sig <= '0';
        wait for 60 ns;
        reset_sig <= '1';
        wait for 6 ns;
        reset_sig <= '0';
        wait for 100 ns;
        
        -- Add additional test cases here if needed

        -- End the simulation
        wait;
    end process;
end testbench_architecture;
