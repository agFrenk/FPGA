mopeps@desklukz.1671:1688891080