library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity fusionator is
  generic (
    WIDTH : integer := 128
  );
  port (
    clk           : in std_logic;
    rst             : in std_logic;
    in_ready_1        : in std_logic;
    in_ready_2        : in std_logic;
    input_1         : in std_logic_vector(WIDTH-1 downto 0);  -- primer input
    size_1          : in integer;   -- size del input 1
    input_2         : in std_logic_vector(WIDTH-1 downto 0);  -- segundo input
    size_2          : in integer;   -- size del input 2
    output          : out std_logic_vector((WIDTH*2)-1 downto 0);   -- output
    out_ready       : out std_logic
    );
end entity fusionator;

architecture structural of fusionator is
  signal output_sig : std_logic_vector(output'range) := (others => '0');  -- senial de output
  signal out_ready_sig : std_logic := '0';  -- senial para output ready


begin  -- architecture structural

  process(clk)
    signal first_element_input2 : std_logic_vector(character_index downto 0 ); 
    signal first_element_input2_count : std_logic_vector(character_index downto 0 ); 
    signal last_element_input1 : integer; 
    signal last_element_input1_count  : integer; 
  begin
    if (clk'event and clk = '1' and in_ready_1 = '1' and in_ready_2 = '1') then
      first_element_input2 <= get_character_from_array(input_2, 1, character_size);
      first_element_input2_count <= to_integer(get_character_from_array(input_2, 0, character_size);)
  
      last_element_input1 <= get_character_from_array(input_1, (size_1 - 1), character_size);  -- aca no estoy seguro si va el -1 o no 
      last_element_input1_count <= to_integer(get_character_from_array(input_1, size_1 - 2, character_size);)

      if(first_element_input2 = last_element_input1) then 
      (output_sig(
        (WIDTH*2)-1 downto ((WIDTH*2) - size_1))
       ) <= input_1(WIDTH - 1 downto (WIDTH -size_1));
      
       -- Seteo el ultimo count como la suma
       (output_sig(
        (WIDTH*2) - size_1 - (2*character_size) - 1 downto ((WIDTH*2) - size_1 - character_size))
       ) <= std_logic_vector(to_unsigned(first_element_input2_count + last_element_input1_count , character_size));
      
       -- Escribo 2*character_set menos de el input_2.
       (output_sig(
        (WIDTH*2) - 1 - size_1 downto ((WIDTH*2) - size_1 - size_2 - (2*character_size)))
       ) <= input_2(WIDTH - 1 - (2*character_size) downto (WIDTH - size_2));

      else 
        (output_sig(
          (WIDTH*2)-1 downto ((WIDTH*2) - size_1))
         ) <= input_1(WIDTH - 1 downto (WIDTH -size_1));
        (output_sig(
          (WIDTH*2)-1 - size_1 downto ((WIDTH*2) - size_1 - size_2))
         ) <= input_2(WIDTH - 1 downto (WIDTH - size_2));

      end if; 
      out_ready_sig <= '1';
    end if; 
  end process;

  output <= output_sig;
  out_ready <= out_ready_sig;

end architecture structural;

